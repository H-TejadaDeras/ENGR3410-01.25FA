/*
 * top comment
 */
`begin_keywords "1800-2005" // SystemVerilog-2005

module top(
    input  logic clk,
    output logic RGB_R,
    output logic RGB_G,
    output logic RGB_B
    );
    
    // Net Declarations
    logic 

    initial begin
        pass
    end
endmodule
`end_keywords "1800-2005" // SystemVerilog-2005